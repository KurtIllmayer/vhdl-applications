---------------------------------------------------------------------------------
-- MIT License

-- Copyright (c) 2019 Kurt Illmayer

-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:

-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.

-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
---------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity multiplier is
 PORT(a_i        : IN   std_ulogic_vector(3 DOWNTO 0);
      b_i        : IN   std_ulogic_vector(3 DOWNTO 0);
      result_o   : OUT  std_ulogic_vector(7 DOWNTO 0));
end multiplier;

architecture Behavioral of multiplier is

 signal result_mult : unsigned(7 downto 0);

begin

  result_mult(7 downto 0) <= unsigned(to_stdlogicvector(a_i(3 downto 0))) * unsigned(to_stdlogicvector(b_i(3 downto 0)));

-- result_o(7 downto 0) <= to_stdulogicvector(result_mult(7 downto 0));
 
--  result_o(7 downto 0) <= to_stdulogicvector(unsigned(to_stdlogicvector(a_i(3 downto 0))) * unsigned(to_stdlogicvector(b_i(3 downto 0))));

  result_o(7 downto 0) <= to_stdulogicvector(conv_std_logic_vector(conv_integer(result_mult(7 downto 0)),8));

end Behavioral;
