---------------------------------------------------------------------------------
-- MIT License

-- Copyright (c) 2019 Kurt Illmayer

-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:

-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.

-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
---------------------------------------------------------------------------------

-----------------------------------------------------------------------
-- Please read the following article on the web regarding the
-- vga video timings:
-- http://www.epanorama.net/documents/pc/vga_timing.html
--
-- This module generates the video synch pulses for the monitor to
-- enter 640x480@60Hz resolution state. The video_enable_o
-- signal is active, when the pixel is inside the visible screen.
-- The color red_o, green_o and blue_o outputs should be reset to 0,
-- when the pixel is outside the visible screen.

-- Timing diagram for the horizontal synch signal (h_sync_o)
-- 0                  640  656    752             799 (pixels)
-- -------------------------|______|-----------------

-- Timing diagram for the vertical synch signal (v_sync_o)
-- 0                            480  490    492   524 (lines)
-- -----------------------------------|______|-------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity vga_controller is
port(-- 100 MHz clock fecg external quartz oscillator
     clk_i          : in  std_ulogic; 
     -- System Reset Signal
     reset_i        : in  std_ulogic; 
      -- Horizontal sync pulse
     h_sync_o       : out std_ulogic; 
     -- Vertical sync pulse   
     v_sync_o       : out std_ulogic;
     -- Output signal for color red
     red_o          : out std_ulogic_vector(2 downto 0); 
     -- Output signal for color green
     green_o        : out std_ulogic_vector(2 downto 0);
     -- Output signal for color blue
     blue_o         : out std_ulogic_vector(1 downto 0));
end vga_controller;

architecture Behavioral of vga_controller is
 -- image clock
 signal clk_25MHz           : std_ulogic;
 -- counter for clock divider
 signal counter             : integer range 0 to 1;
 -- signal for coclor red
 signal red, red_blacked    : std_ulogic_vector(2 downto 0);
 -- signal for coclor green
 signal green, green_blacked: std_ulogic_vector(2 downto 0);
 -- signal for color blue
 signal blue, blue_blacked  : std_ulogic_vector(1 downto 0);
 -- maximum value for the horizontal pixel counter
 constant h_max_c           : std_logic_vector(9 downto 0) := "1100100000"; -- 800
 -- maximum value for the vertical pixel counter
 constant v_max_c           : std_logic_vector(9 downto 0) := "1000001101"; -- 525
 -- total number of visible columns
 constant h_pixels_c        : std_logic_vector(9 downto 0) := "1010000000"; -- 640
 -- value for the horizontal counter where front porch ends
 constant h_front_porch_c   : std_logic_vector(9 downto 0) := "1010010000"; -- 656
 -- value for the horizontal counter where the synch pulse ends
 constant h_sync_pulse_c    : std_logic_vector(9 downto 0) := "1011110000"; -- 752
 -- total number of visible lines
 constant v_lines_c         : std_logic_vector(9 downto 0) := "0111100000"; -- 480
 -- total number of visible lines
 constant v_distance_c      : std_logic_vector(9 downto 0) := "0100101100"; -- 300 
 -- value for the vertical counter where the front porch ends
 constant v_front_porch_c   : std_logic_vector(9 downto 0) := "0111101010"; -- 490
 -- value for the vertical counter where the synch pulse ends
 constant v_sync_pulse_c    : std_logic_vector(9 downto 0) := "0111101100"; -- 492
 -- horizontal counter
 signal h_counter           : std_logic_vector(9 downto 0);
 -- vertical counter
 signal v_counter           : std_logic_vector(9 downto 0);
 -- enables the three colors: red, green and blue
 signal video_enable        : std_ulogic;
 -- clock for blacked video lines
 signal clk_64Hz            : std_ulogic; 
 -- clock divider for clk_64Hz
 signal counter_64          : integer range 0 to 781249;
 -- Count signal for black signal: 10 x signal with 64 pixels
 signal count_black         : integer range 0 to 639;   
 -- Maximum count value for black signal
 constant count_max_c       : integer range 0 to 639 := 639;
 -- Data from the ecg diagram
 type rom_640 is array (0 to 639) of std_logic_vector(5 downto 0);
  
   -------------------------------------------------------------------------------  
   -- Put here your ECG Curve with 64 vaues 10 times one after another:
   -- So you get 64*10 = 640 values:
   -------------------------------------------------------------------------------   
   constant ecg : rom_640 :=
	("000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
    "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
    "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
    "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000111",
	 "001001",
	 "001011",
	 "001110",
	 "010000",
	 "010001",
	 "010000",
	 "001110",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
 	 "000110",
	 "000010",
	 "000110",
	 "010010",
	 "100100",
	 "101101",
	 "110111",
	 "111111",
	 "110111",
	 "101101",
	 "100100",
	 "010010",
	 "000110",
	 "000000",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "001001",
	 "001011",
	 "001111",
	 "010011",
	 "010110",
	 "010111",
	 "010110",
	 "010011",
	 "001111",
	 "001011",
	 "001001",
	 "000111",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110",
	 "000110");    
   -------------------------------------------------------------------------------

begin

   -- clock_divider   
   divide_p: process(clk_i, reset_i)
   begin   
      if(reset_i = '1')then
          counter   <=  0;
          clk_25MHz <= '0';          
      elsif(clk_i'event and clk_i ='1') then
         if(counter = 1) then
            counter   <= 0;
            clk_25MHz <= not clk_25MHz;
         else
            counter   <= counter + 1;
         end if;
      end if;
   end process divide_p;

   -- increment horizontal counter at clk_25MHz rate
   -- until h_max_c is reached, then reset and keep counting
   h_count_p: process(clk_25MHz, reset_i)
   begin   
      if(reset_i = '1')then
          h_counter <= (others => '0');      
      elsif(clk_25MHz'event and clk_25MHz ='1') then
         if(h_counter = h_max_c - "0000000001") then
            h_counter <= (others => '0');
         else
            h_counter <= h_counter + "0000000001";
         end if;
      end if;
   end process h_count_p;

   -- increment vertical counter when one line is finished
   -- (horizontal counter reached h_max_c)
   -- until v_max_c is reached, then reset and keep counting
   v_count_p: process(clk_25MHz, reset_i)
   begin
      if(reset_i = '1')then
          v_counter <= (others => '0');     
      elsif(clk_25MHz'event and clk_25MHz ='1') then
         if(h_counter = h_max_c - "0000000001") then
            if(v_counter = v_max_c - "0000000001") then
               v_counter <= (others => '0');
            else
               v_counter <= v_counter + "0000000001";
            end if;
         end if;
      end if;
   end process v_count_p;

   -- generate horizontal synch pulse when horizontal counter 
   -- is between where the front porch ends and the synch pulse ends.
   -- The h_sync_ois active (with polarity sync_pulse_polarity_c) 
   -- for a total of 96 pixels.
   hs_p: process(clk_25MHz, reset_i)
   begin
      if(reset_i = '1')then
          h_sync_o <= '1';  
      elsif(clk_25MHz'event and clk_25MHz ='1') then
         if((h_counter >= h_front_porch_c) and (h_counter < h_sync_pulse_c)) then
            h_sync_o <= '0';
         else
            h_sync_o <= '1';
         end if;
      end if;
   end process hs_p;

   -- generate vertical synch pulse
   -- when vertical counter is between where the
   -- front porch ends and the synch pulse ends.
   -- The v_sync_ois active (with polarity sync_pulse_polarity_c) 
   -- for a total of 2 video lines = 2*h_max_c = 1600 pixels.
   vs_p: process(clk_25MHz, reset_i)
   begin
      if(reset_i = '1')then
          v_sync_o <= '1'; 
      elsif(clk_25MHz'event and clk_25MHz ='1') then
         if((v_counter >= v_front_porch_c) and (v_counter < v_sync_pulse_c)) then
            v_sync_o <= '0';
         else
            v_sync_o <= '1';
         end if;
      end if;
   end process vs_p;

   --  enable video output when pixel is in visible area
   video_p: process(clk_25MHz, reset_i)
   begin
      if(reset_i = '1')then
          video_enable <= '0';       
      elsif(clk_25MHz'event and clk_25MHz ='1') then
         -- Visible image range
         if((h_counter < h_pixels_c) and (v_counter < v_lines_c)) then
            video_enable <= '1';
         else
            video_enable <= '0';
         end if;
      end if;
   end process video_p;
 
   red_o   <=   red_blacked when video_enable = '1' else "000";

   green_o <= green_blacked when video_enable = '1' else "000";

   blue_o  <=  blue_blacked when video_enable = '1' else  "00";
 
   divide_64_p: process(clk_i, reset_i)
   begin   
      if(reset_i = '1')then
          counter_64   <=  0;
          clk_64Hz     <= '0';          
      elsif(clk_i'event and clk_i ='1') then
         if(counter_64 = 781249) then
            counter_64   <= 0;
            clk_64Hz     <= not clk_64Hz;
         else
            counter_64   <= counter_64 + 1;
         end if;
      end if;
   end process divide_64_p;
 
   black_p:process(reset_i, clk_64Hz)
   begin
   if(reset_i = '1')then
       count_black <= 0;       
   elsif(clk_64Hz'event and clk_64Hz ='1') then
     if(count_black = count_max_c)then
        count_black <= 0;
     else
        count_black <= count_black + 1;         
     end if;
   end if;     
   end process black_p;   
   
   blacked_p: process(h_counter, count_black, red, green, blue)
   begin                              
   if((h_counter = count_black) or (h_counter = (count_black + 1)) or (h_counter = (count_black + 2))
   or (h_counter = (count_black + 3)) or (h_counter = (count_black + 4)) or (h_counter = (count_black + 5)))then
      red_blacked   <= "000";
      green_blacked <= "000";
      blue_blacked  <=  "00";  
   else
      red_blacked   <=   red;
      green_blacked <= green;
      blue_blacked  <=  blue; 
   end if;
   end process blacked_p;   
  
 image_p: process(reset_i, clk_25MHz, h_counter, v_counter)
 begin                              
                   
 if(reset_i = '1')then
     red   <= "000";
     green <= "000";
     blue  <=  "00";  
 elsif(clk_25MHz'event and clk_25MHz ='1') then
                   
 case h_counter is                    

 when "0000000000" => if(ecg(1) > ecg(0))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(1))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(0)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(1) < ecg(0))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(0))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(1)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(0))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000001" => if(ecg(2) > ecg(1))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(2))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(1)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(2) < ecg(1))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(1))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(2)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(1))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000010" => if(ecg(3) > ecg(2))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(3))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(2)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(3) < ecg(2))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(2))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(3)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(2))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000011" => if(ecg(4) > ecg(3))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(4))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(3)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(4) < ecg(3))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(3))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(4)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(3))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000100" => if(ecg(5) > ecg(4))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(5))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(4)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(5) < ecg(4))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(4))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(5)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(4))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000101" => if(ecg(6) > ecg(5))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(6))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(5)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(6) < ecg(5))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(5))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(6)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(5))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000110" => if(ecg(7) > ecg(6))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(7))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(6)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(7) < ecg(6))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(6))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(7)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(6))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000000111" => if(ecg(8) > ecg(7))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(8))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(7)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(8) < ecg(7))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(7))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(8)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(7))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001000" => if(ecg(9) > ecg(8))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(9))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(8)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(9) < ecg(8))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(8))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(9)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(8))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001001" => if(ecg(10) > ecg(9))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(10))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(9)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(10) < ecg(9))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(9))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(10)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(9))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001010" => if(ecg(11) > ecg(10))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(11))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(10)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(11) < ecg(10))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(10))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(11)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(10))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001011" => if(ecg(12) > ecg(11))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(12))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(11)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(12) < ecg(11))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(11))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(12)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(11))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001100" => if(ecg(13) > ecg(12))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(13))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(12)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(13) < ecg(12))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(12))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(13)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(12))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001101" => if(ecg(14) > ecg(13))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(14))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(13)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(14) < ecg(13))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(13))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(14)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(13))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001110" => if(ecg(15) > ecg(14))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(15))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(14)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(15) < ecg(14))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(14))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(15)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(14))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000001111" => if(ecg(16) > ecg(15))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(16))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(15)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(16) < ecg(15))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(15))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(16)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(15))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010000" => if(ecg(17) > ecg(16))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(17))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(16)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(17) < ecg(16))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(16))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(17)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(16))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010001" => if(ecg(18) > ecg(17))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(18))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(17)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(18) < ecg(17))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(17))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(18)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(17))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010010" => if(ecg(19) > ecg(18))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(19))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(18)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(19) < ecg(18))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(18))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(19)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(18))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010011" => if(ecg(20) > ecg(19))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(20))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(19)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(20) < ecg(19))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(19))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(20)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(19))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010100" => if(ecg(21) > ecg(20))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(21))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(20)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(21) < ecg(20))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(20))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(21)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(20))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010101" => if(ecg(22) > ecg(21))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(22))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(21)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(22) < ecg(21))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(21))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(22)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(21))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010110" => if(ecg(23) > ecg(22))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(23))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(22)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(23) < ecg(22))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(22))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(23)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(22))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000010111" => if(ecg(24) > ecg(23))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(24))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(23)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(24) < ecg(23))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(23))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(24)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(23))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011000" => if(ecg(25) > ecg(24))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(25))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(24)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(25) < ecg(24))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(24))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(25)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(24))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011001" => if(ecg(26) > ecg(25))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(26))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(25)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(26) < ecg(25))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(25))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(26)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(25))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011010" => if(ecg(27) > ecg(26))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(27))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(26)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(27) < ecg(26))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(26))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(27)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(26))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011011" => if(ecg(28) > ecg(27))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(28))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(27)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(28) < ecg(27))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(27))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(28)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(27))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011100" => if(ecg(29) > ecg(28))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(29))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(28)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(29) < ecg(28))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(28))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(29)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(28))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011101" => if(ecg(30) > ecg(29))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(30))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(29)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(30) < ecg(29))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(29))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(30)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(29))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011110" => if(ecg(31) > ecg(30))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(31))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(30)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(31) < ecg(30))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(30))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(31)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(30))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000011111" => if(ecg(32) > ecg(31))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(32))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(31)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(32) < ecg(31))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(31))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(32)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(31))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100000" => if(ecg(33) > ecg(32))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(33))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(32)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(33) < ecg(32))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(32))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(33)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(32))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100001" => if(ecg(34) > ecg(33))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(34))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(33)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(34) < ecg(33))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(33))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(34)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(33))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100010" => if(ecg(35) > ecg(34))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(35))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(34)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(35) < ecg(34))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(34))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(35)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(34))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100011" => if(ecg(36) > ecg(35))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(36))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(35)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(36) < ecg(35))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(35))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(36)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(35))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100100" => if(ecg(37) > ecg(36))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(37))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(36)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(37) < ecg(36))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(36))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(37)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(36))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100101" => if(ecg(38) > ecg(37))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(38))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(37)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(38) < ecg(37))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(37))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(38)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(37))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100110" => if(ecg(39) > ecg(38))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(39))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(38)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(39) < ecg(38))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(38))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(39)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(38))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000100111" => if(ecg(40) > ecg(39))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(40))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(39)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(40) < ecg(39))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(39))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(40)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(39))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101000" => if(ecg(41) > ecg(40))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(41))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(40)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(41) < ecg(40))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(40))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(41)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(40))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101001" => if(ecg(42) > ecg(41))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(42))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(41)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(42) < ecg(41))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(41))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(42)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(41))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101010" => if(ecg(43) > ecg(42))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(43))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(42)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(43) < ecg(42))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(42))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(43)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(42))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101011" => if(ecg(44) > ecg(43))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(44))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(43)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(44) < ecg(43))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(43))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(44)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(43))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101100" => if(ecg(45) > ecg(44))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(45))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(44)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(45) < ecg(44))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(44))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(45)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(44))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101101" => if(ecg(46) > ecg(45))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(46))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(45)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(46) < ecg(45))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(45))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(46)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(45))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101110" => if(ecg(47) > ecg(46))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(47))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(46)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(47) < ecg(46))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(46))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(47)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(46))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000101111" => if(ecg(48) > ecg(47))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(48))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(47)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(48) < ecg(47))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(47))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(48)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(47))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110000" => if(ecg(49) > ecg(48))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(49))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(48)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(49) < ecg(48))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(48))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(49)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(48))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110001" => if(ecg(50) > ecg(49))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(50))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(49)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(50) < ecg(49))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(49))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(50)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(49))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110010" => if(ecg(51) > ecg(50))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(51))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(50)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(51) < ecg(50))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(50))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(51)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(50))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110011" => if(ecg(52) > ecg(51))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(52))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(51)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(52) < ecg(51))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(51))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(52)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(51))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110100" => if(ecg(53) > ecg(52))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(53))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(52)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(53) < ecg(52))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(52))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(53)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(52))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110101" => if(ecg(54) > ecg(53))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(54))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(53)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(54) < ecg(53))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(53))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(54)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(53))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110110" => if(ecg(55) > ecg(54))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(55))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(54)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(55) < ecg(54))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(54))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(55)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(54))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000110111" => if(ecg(56) > ecg(55))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(56))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(55)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(56) < ecg(55))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(55))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(56)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(55))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111000" => if(ecg(57) > ecg(56))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(57))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(56)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(57) < ecg(56))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(56))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(57)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(56))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111001" => if(ecg(58) > ecg(57))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(58))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(57)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(58) < ecg(57))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(57))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(58)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(57))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111010" => if(ecg(59) > ecg(58))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(59))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(58)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(59) < ecg(58))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(58))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(59)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(58))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111011" => if(ecg(60) > ecg(59))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(60))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(59)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(60) < ecg(59))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(59))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(60)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(59))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111100" => if(ecg(61) > ecg(60))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(61))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(60)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(61) < ecg(60))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(60))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(61)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(60))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111101" => if(ecg(62) > ecg(61))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(62))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(61)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(62) < ecg(61))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(61))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(62)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(61))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111110" => if(ecg(63) > ecg(62))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(63))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(62)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(63) < ecg(62))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(62))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(63)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(62))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0000111111" => if(ecg(64) > ecg(63))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(64))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(63)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(64) < ecg(63))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(63))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(64)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(63))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000000" => if(ecg(65) > ecg(64))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(65))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(64)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(65) < ecg(64))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(64))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(65)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(64))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000001" => if(ecg(66) > ecg(65))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(66))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(65)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(66) < ecg(65))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(65))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(66)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(65))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000010" => if(ecg(67) > ecg(66))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(67))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(66)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(67) < ecg(66))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(66))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(67)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(66))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000011" => if(ecg(68) > ecg(67))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(68))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(67)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(68) < ecg(67))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(67))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(68)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(67))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000100" => if(ecg(69) > ecg(68))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(69))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(68)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(69) < ecg(68))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(68))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(69)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(68))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000101" => if(ecg(70) > ecg(69))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(70))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(69)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(70) < ecg(69))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(69))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(70)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(69))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000110" => if(ecg(71) > ecg(70))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(71))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(70)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(71) < ecg(70))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(70))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(71)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(70))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001000111" => if(ecg(72) > ecg(71))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(72))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(71)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(72) < ecg(71))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(71))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(72)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(71))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001000" => if(ecg(73) > ecg(72))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(73))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(72)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(73) < ecg(72))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(72))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(73)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(72))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001001" => if(ecg(74) > ecg(73))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(74))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(73)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(74) < ecg(73))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(73))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(74)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(73))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001010" => if(ecg(75) > ecg(74))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(75))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(74)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(75) < ecg(74))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(74))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(75)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(74))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001011" => if(ecg(76) > ecg(75))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(76))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(75)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(76) < ecg(75))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(75))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(76)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(75))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001100" => if(ecg(77) > ecg(76))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(77))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(76)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(77) < ecg(76))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(76))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(77)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(76))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001101" => if(ecg(78) > ecg(77))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(78))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(77)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(78) < ecg(77))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(77))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(78)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(77))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001110" => if(ecg(79) > ecg(78))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(79))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(78)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(79) < ecg(78))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(78))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(79)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(78))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001001111" => if(ecg(80) > ecg(79))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(80))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(79)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(80) < ecg(79))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(79))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(80)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(79))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010000" => if(ecg(81) > ecg(80))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(81))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(80)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(81) < ecg(80))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(80))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(81)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(80))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010001" => if(ecg(82) > ecg(81))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(82))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(81)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(82) < ecg(81))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(81))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(82)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(81))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010010" => if(ecg(83) > ecg(82))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(83))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(82)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(83) < ecg(82))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(82))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(83)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(82))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010011" => if(ecg(84) > ecg(83))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(84))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(83)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(84) < ecg(83))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(83))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(84)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(83))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010100" => if(ecg(85) > ecg(84))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(85))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(84)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(85) < ecg(84))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(84))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(85)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(84))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010101" => if(ecg(86) > ecg(85))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(86))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(85)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(86) < ecg(85))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(85))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(86)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(85))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010110" => if(ecg(87) > ecg(86))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(87))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(86)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(87) < ecg(86))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(86))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(87)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(86))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001010111" => if(ecg(88) > ecg(87))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(88))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(87)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(88) < ecg(87))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(87))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(88)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(87))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011000" => if(ecg(89) > ecg(88))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(89))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(88)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(89) < ecg(88))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(88))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(89)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(88))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011001" => if(ecg(90) > ecg(89))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(90))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(89)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(90) < ecg(89))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(89))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(90)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(89))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011010" => if(ecg(91) > ecg(90))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(91))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(90)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(91) < ecg(90))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(90))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(91)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(90))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011011" => if(ecg(92) > ecg(91))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(92))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(91)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(92) < ecg(91))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(91))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(92)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(91))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011100" => if(ecg(93) > ecg(92))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(93))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(92)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(93) < ecg(92))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(92))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(93)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(92))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011101" => if(ecg(94) > ecg(93))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(94))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(93)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(94) < ecg(93))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(93))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(94)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(93))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011110" => if(ecg(95) > ecg(94))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(95))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(94)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(95) < ecg(94))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(94))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(95)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(94))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001011111" => if(ecg(96) > ecg(95))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(96))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(95)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(96) < ecg(95))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(95))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(96)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(95))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100000" => if(ecg(97) > ecg(96))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(97))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(96)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(97) < ecg(96))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(96))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(97)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(96))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100001" => if(ecg(98) > ecg(97))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(98))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(97)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(98) < ecg(97))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(97))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(98)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(97))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100010" => if(ecg(99) > ecg(98))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(99))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(98)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(99) < ecg(98))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(98))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(99)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(98))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100011" => if(ecg(100) > ecg(99))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(100))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(99)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(100) < ecg(99))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(99))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(100)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(99))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100100" => if(ecg(101) > ecg(100))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(101))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(100)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(101) < ecg(100))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(100))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(101)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(100))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100101" => if(ecg(102) > ecg(101))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(102))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(101)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(102) < ecg(101))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(101))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(102)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(101))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100110" => if(ecg(103) > ecg(102))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(103))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(102)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(103) < ecg(102))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(102))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(103)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(102))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001100111" => if(ecg(104) > ecg(103))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(104))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(103)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(104) < ecg(103))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(103))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(104)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(103))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101000" => if(ecg(105) > ecg(104))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(105))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(104)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(105) < ecg(104))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(104))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(105)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(104))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101001" => if(ecg(106) > ecg(105))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(106))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(105)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(106) < ecg(105))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(105))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(106)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(105))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101010" => if(ecg(107) > ecg(106))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(107))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(106)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(107) < ecg(106))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(106))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(107)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(106))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101011" => if(ecg(108) > ecg(107))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(108))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(107)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(108) < ecg(107))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(107))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(108)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(107))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101100" => if(ecg(109) > ecg(108))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(109))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(108)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(109) < ecg(108))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(108))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(109)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(108))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101101" => if(ecg(110) > ecg(109))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(110))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(109)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(110) < ecg(109))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(109))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(110)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(109))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101110" => if(ecg(111) > ecg(110))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(111))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(110)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(111) < ecg(110))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(110))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(111)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(110))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001101111" => if(ecg(112) > ecg(111))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(112))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(111)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(112) < ecg(111))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(111))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(112)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(111))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110000" => if(ecg(113) > ecg(112))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(113))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(112)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(113) < ecg(112))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(112))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(113)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(112))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110001" => if(ecg(114) > ecg(113))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(114))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(113)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(114) < ecg(113))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(113))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(114)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(113))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110010" => if(ecg(115) > ecg(114))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(115))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(114)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(115) < ecg(114))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(114))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(115)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(114))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110011" => if(ecg(116) > ecg(115))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(116))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(115)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(116) < ecg(115))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(115))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(116)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(115))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110100" => if(ecg(117) > ecg(116))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(117))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(116)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(117) < ecg(116))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(116))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(117)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(116))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110101" => if(ecg(118) > ecg(117))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(118))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(117)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(118) < ecg(117))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(117))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(118)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(117))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110110" => if(ecg(119) > ecg(118))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(119))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(118)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(119) < ecg(118))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(118))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(119)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(118))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001110111" => if(ecg(120) > ecg(119))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(120))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(119)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(120) < ecg(119))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(119))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(120)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(119))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111000" => if(ecg(121) > ecg(120))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(121))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(120)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(121) < ecg(120))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(120))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(121)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(120))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111001" => if(ecg(122) > ecg(121))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(122))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(121)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(122) < ecg(121))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(121))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(122)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(121))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111010" => if(ecg(123) > ecg(122))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(123))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(122)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(123) < ecg(122))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(122))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(123)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(122))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111011" => if(ecg(124) > ecg(123))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(124))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(123)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(124) < ecg(123))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(123))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(124)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(123))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111100" => if(ecg(125) > ecg(124))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(125))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(124)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(125) < ecg(124))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(124))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(125)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(124))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111101" => if(ecg(126) > ecg(125))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(126))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(125)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(126) < ecg(125))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(125))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(126)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(125))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111110" => if(ecg(127) > ecg(126))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(127))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(126)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(127) < ecg(126))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(126))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(127)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(126))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0001111111" => if(ecg(128) > ecg(127))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(128))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(127)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(128) < ecg(127))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(127))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(128)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(127))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000000" => if(ecg(129) > ecg(128))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(129))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(128)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(129) < ecg(128))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(128))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(129)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(128))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000001" => if(ecg(130) > ecg(129))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(130))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(129)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(130) < ecg(129))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(129))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(130)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(129))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000010" => if(ecg(131) > ecg(130))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(131))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(130)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(131) < ecg(130))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(130))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(131)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(130))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000011" => if(ecg(132) > ecg(131))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(132))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(131)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(132) < ecg(131))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(131))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(132)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(131))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000100" => if(ecg(133) > ecg(132))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(133))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(132)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(133) < ecg(132))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(132))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(133)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(132))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000101" => if(ecg(134) > ecg(133))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(134))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(133)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(134) < ecg(133))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(133))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(134)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(133))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000110" => if(ecg(135) > ecg(134))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(135))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(134)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(135) < ecg(134))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(134))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(135)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(134))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010000111" => if(ecg(136) > ecg(135))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(136))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(135)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(136) < ecg(135))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(135))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(136)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(135))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001000" => if(ecg(137) > ecg(136))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(137))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(136)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(137) < ecg(136))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(136))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(137)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(136))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001001" => if(ecg(138) > ecg(137))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(138))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(137)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(138) < ecg(137))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(137))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(138)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(137))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001010" => if(ecg(139) > ecg(138))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(139))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(138)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(139) < ecg(138))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(138))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(139)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(138))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001011" => if(ecg(140) > ecg(139))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(140))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(139)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(140) < ecg(139))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(139))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(140)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(139))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001100" => if(ecg(141) > ecg(140))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(141))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(140)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(141) < ecg(140))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(140))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(141)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(140))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001101" => if(ecg(142) > ecg(141))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(142))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(141)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(142) < ecg(141))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(141))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(142)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(141))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001110" => if(ecg(143) > ecg(142))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(143))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(142)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(143) < ecg(142))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(142))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(143)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(142))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010001111" => if(ecg(144) > ecg(143))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(144))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(143)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(144) < ecg(143))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(143))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(144)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(143))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010000" => if(ecg(145) > ecg(144))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(145))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(144)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(145) < ecg(144))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(144))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(145)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(144))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010001" => if(ecg(146) > ecg(145))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(146))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(145)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(146) < ecg(145))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(145))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(146)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(145))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010010" => if(ecg(147) > ecg(146))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(147))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(146)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(147) < ecg(146))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(146))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(147)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(146))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010011" => if(ecg(148) > ecg(147))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(148))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(147)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(148) < ecg(147))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(147))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(148)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(147))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010100" => if(ecg(149) > ecg(148))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(149))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(148)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(149) < ecg(148))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(148))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(149)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(148))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010101" => if(ecg(150) > ecg(149))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(150))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(149)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(150) < ecg(149))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(149))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(150)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(149))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010110" => if(ecg(151) > ecg(150))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(151))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(150)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(151) < ecg(150))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(150))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(151)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(150))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010010111" => if(ecg(152) > ecg(151))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(152))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(151)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(152) < ecg(151))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(151))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(152)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(151))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011000" => if(ecg(153) > ecg(152))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(153))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(152)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(153) < ecg(152))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(152))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(153)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(152))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011001" => if(ecg(154) > ecg(153))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(154))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(153)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(154) < ecg(153))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(153))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(154)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(153))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011010" => if(ecg(155) > ecg(154))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(155))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(154)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(155) < ecg(154))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(154))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(155)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(154))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011011" => if(ecg(156) > ecg(155))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(156))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(155)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(156) < ecg(155))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(155))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(156)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(155))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011100" => if(ecg(157) > ecg(156))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(157))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(156)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(157) < ecg(156))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(156))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(157)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(156))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011101" => if(ecg(158) > ecg(157))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(158))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(157)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(158) < ecg(157))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(157))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(158)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(157))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011110" => if(ecg(159) > ecg(158))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(159))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(158)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(159) < ecg(158))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(158))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(159)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(158))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010011111" => if(ecg(160) > ecg(159))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(160))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(159)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(160) < ecg(159))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(159))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(160)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(159))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100000" => if(ecg(161) > ecg(160))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(161))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(160)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(161) < ecg(160))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(160))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(161)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(160))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100001" => if(ecg(162) > ecg(161))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(162))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(161)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(162) < ecg(161))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(161))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(162)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(161))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100010" => if(ecg(163) > ecg(162))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(163))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(162)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(163) < ecg(162))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(162))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(163)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(162))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100011" => if(ecg(164) > ecg(163))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(164))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(163)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(164) < ecg(163))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(163))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(164)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(163))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100100" => if(ecg(165) > ecg(164))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(165))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(164)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(165) < ecg(164))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(164))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(165)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(164))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100101" => if(ecg(166) > ecg(165))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(166))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(165)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(166) < ecg(165))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(165))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(166)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(165))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100110" => if(ecg(167) > ecg(166))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(167))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(166)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(167) < ecg(166))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(166))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(167)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(166))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010100111" => if(ecg(168) > ecg(167))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(168))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(167)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(168) < ecg(167))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(167))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(168)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(167))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101000" => if(ecg(169) > ecg(168))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(169))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(168)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(169) < ecg(168))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(168))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(169)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(168))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101001" => if(ecg(170) > ecg(169))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(170))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(169)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(170) < ecg(169))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(169))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(170)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(169))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101010" => if(ecg(171) > ecg(170))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(171))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(170)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(171) < ecg(170))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(170))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(171)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(170))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101011" => if(ecg(172) > ecg(171))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(172))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(171)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(172) < ecg(171))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(171))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(172)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(171))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101100" => if(ecg(173) > ecg(172))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(173))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(172)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(173) < ecg(172))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(172))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(173)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(172))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101101" => if(ecg(174) > ecg(173))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(174))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(173)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(174) < ecg(173))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(173))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(174)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(173))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101110" => if(ecg(175) > ecg(174))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(175))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(174)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(175) < ecg(174))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(174))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(175)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(174))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010101111" => if(ecg(176) > ecg(175))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(176))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(175)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(176) < ecg(175))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(175))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(176)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(175))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110000" => if(ecg(177) > ecg(176))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(177))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(176)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(177) < ecg(176))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(176))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(177)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(176))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110001" => if(ecg(178) > ecg(177))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(178))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(177)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(178) < ecg(177))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(177))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(178)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(177))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110010" => if(ecg(179) > ecg(178))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(179))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(178)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(179) < ecg(178))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(178))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(179)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(178))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110011" => if(ecg(180) > ecg(179))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(180))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(179)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(180) < ecg(179))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(179))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(180)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(179))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110100" => if(ecg(181) > ecg(180))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(181))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(180)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(181) < ecg(180))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(180))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(181)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(180))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110101" => if(ecg(182) > ecg(181))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(182))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(181)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(182) < ecg(181))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(181))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(182)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(181))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110110" => if(ecg(183) > ecg(182))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(183))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(182)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(183) < ecg(182))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(182))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(183)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(182))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010110111" => if(ecg(184) > ecg(183))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(184))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(183)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(184) < ecg(183))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(183))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(184)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(183))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111000" => if(ecg(185) > ecg(184))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(185))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(184)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(185) < ecg(184))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(184))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(185)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(184))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111001" => if(ecg(186) > ecg(185))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(186))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(185)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(186) < ecg(185))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(185))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(186)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(185))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111010" => if(ecg(187) > ecg(186))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(187))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(186)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(187) < ecg(186))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(186))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(187)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(186))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111011" => if(ecg(188) > ecg(187))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(188))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(187)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(188) < ecg(187))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(187))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(188)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(187))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111100" => if(ecg(189) > ecg(188))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(189))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(188)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(189) < ecg(188))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(188))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(189)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(188))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111101" => if(ecg(190) > ecg(189))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(190))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(189)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(190) < ecg(189))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(189))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(190)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(189))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111110" => if(ecg(191) > ecg(190))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(191))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(190)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(191) < ecg(190))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(190))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(191)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(190))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0010111111" => if(ecg(192) > ecg(191))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(192))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(191)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(192) < ecg(191))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(191))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(192)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(191))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000000" => if(ecg(193) > ecg(192))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(193))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(192)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(193) < ecg(192))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(192))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(193)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(192))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000001" => if(ecg(194) > ecg(193))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(194))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(193)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(194) < ecg(193))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(193))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(194)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(193))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000010" => if(ecg(195) > ecg(194))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(195))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(194)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(195) < ecg(194))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(194))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(195)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(194))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000011" => if(ecg(196) > ecg(195))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(196))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(195)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(196) < ecg(195))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(195))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(196)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(195))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000100" => if(ecg(197) > ecg(196))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(197))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(196)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(197) < ecg(196))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(196))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(197)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(196))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000101" => if(ecg(198) > ecg(197))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(198))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(197)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(198) < ecg(197))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(197))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(198)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(197))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000110" => if(ecg(199) > ecg(198))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(199))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(198)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(199) < ecg(198))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(198))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(199)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(198))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011000111" => if(ecg(200) > ecg(199))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(200))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(199)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(200) < ecg(199))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(199))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(200)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(199))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001000" => if(ecg(201) > ecg(200))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(201))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(200)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(201) < ecg(200))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(200))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(201)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(200))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001001" => if(ecg(202) > ecg(201))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(202))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(201)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(202) < ecg(201))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(201))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(202)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(201))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001010" => if(ecg(203) > ecg(202))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(203))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(202)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(203) < ecg(202))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(202))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(203)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(202))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001011" => if(ecg(204) > ecg(203))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(204))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(203)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(204) < ecg(203))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(203))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(204)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(203))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001100" => if(ecg(205) > ecg(204))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(205))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(204)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(205) < ecg(204))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(204))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(205)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(204))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001101" => if(ecg(206) > ecg(205))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(206))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(205)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(206) < ecg(205))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(205))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(206)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(205))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001110" => if(ecg(207) > ecg(206))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(207))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(206)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(207) < ecg(206))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(206))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(207)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(206))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011001111" => if(ecg(208) > ecg(207))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(208))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(207)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(208) < ecg(207))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(207))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(208)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(207))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010000" => if(ecg(209) > ecg(208))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(209))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(208)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(209) < ecg(208))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(208))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(209)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(208))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010001" => if(ecg(210) > ecg(209))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(210))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(209)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(210) < ecg(209))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(209))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(210)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(209))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010010" => if(ecg(211) > ecg(210))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(211))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(210)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(211) < ecg(210))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(210))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(211)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(210))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010011" => if(ecg(212) > ecg(211))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(212))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(211)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(212) < ecg(211))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(211))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(212)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(211))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010100" => if(ecg(213) > ecg(212))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(213))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(212)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(213) < ecg(212))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(212))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(213)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(212))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010101" => if(ecg(214) > ecg(213))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(214))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(213)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(214) < ecg(213))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(213))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(214)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(213))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010110" => if(ecg(215) > ecg(214))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(215))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(214)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(215) < ecg(214))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(214))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(215)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(214))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011010111" => if(ecg(216) > ecg(215))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(216))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(215)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(216) < ecg(215))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(215))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(216)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(215))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011000" => if(ecg(217) > ecg(216))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(217))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(216)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(217) < ecg(216))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(216))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(217)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(216))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011001" => if(ecg(218) > ecg(217))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(218))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(217)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(218) < ecg(217))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(217))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(218)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(217))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011010" => if(ecg(219) > ecg(218))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(219))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(218)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(219) < ecg(218))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(218))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(219)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(218))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011011" => if(ecg(220) > ecg(219))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(220))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(219)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(220) < ecg(219))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(219))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(220)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(219))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011100" => if(ecg(221) > ecg(220))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(221))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(220)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(221) < ecg(220))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(220))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(221)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(220))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011101" => if(ecg(222) > ecg(221))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(222))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(221)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(222) < ecg(221))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(221))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(222)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(221))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011110" => if(ecg(223) > ecg(222))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(223))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(222)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(223) < ecg(222))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(222))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(223)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(222))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011011111" => if(ecg(224) > ecg(223))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(224))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(223)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(224) < ecg(223))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(223))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(224)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(223))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100000" => if(ecg(225) > ecg(224))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(225))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(224)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(225) < ecg(224))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(224))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(225)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(224))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100001" => if(ecg(226) > ecg(225))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(226))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(225)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(226) < ecg(225))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(225))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(226)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(225))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100010" => if(ecg(227) > ecg(226))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(227))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(226)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(227) < ecg(226))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(226))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(227)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(226))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100011" => if(ecg(228) > ecg(227))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(228))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(227)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(228) < ecg(227))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(227))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(228)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(227))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100100" => if(ecg(229) > ecg(228))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(229))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(228)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(229) < ecg(228))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(228))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(229)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(228))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100101" => if(ecg(230) > ecg(229))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(230))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(229)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(230) < ecg(229))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(229))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(230)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(229))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100110" => if(ecg(231) > ecg(230))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(231))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(230)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(231) < ecg(230))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(230))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(231)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(230))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011100111" => if(ecg(232) > ecg(231))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(232))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(231)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(232) < ecg(231))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(231))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(232)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(231))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101000" => if(ecg(233) > ecg(232))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(233))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(232)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(233) < ecg(232))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(232))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(233)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(232))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101001" => if(ecg(234) > ecg(233))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(234))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(233)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(234) < ecg(233))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(233))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(234)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(233))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101010" => if(ecg(235) > ecg(234))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(235))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(234)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(235) < ecg(234))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(234))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(235)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(234))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101011" => if(ecg(236) > ecg(235))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(236))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(235)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(236) < ecg(235))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(235))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(236)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(235))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101100" => if(ecg(237) > ecg(236))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(237))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(236)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(237) < ecg(236))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(236))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(237)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(236))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101101" => if(ecg(238) > ecg(237))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(238))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(237)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(238) < ecg(237))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(237))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(238)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(237))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101110" => if(ecg(239) > ecg(238))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(239))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(238)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(239) < ecg(238))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(238))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(239)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(238))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011101111" => if(ecg(240) > ecg(239))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(240))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(239)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(240) < ecg(239))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(239))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(240)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(239))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110000" => if(ecg(241) > ecg(240))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(241))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(240)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(241) < ecg(240))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(240))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(241)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(240))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110001" => if(ecg(242) > ecg(241))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(242))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(241)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(242) < ecg(241))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(241))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(242)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(241))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110010" => if(ecg(243) > ecg(242))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(243))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(242)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(243) < ecg(242))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(242))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(243)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(242))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110011" => if(ecg(244) > ecg(243))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(244))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(243)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(244) < ecg(243))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(243))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(244)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(243))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110100" => if(ecg(245) > ecg(244))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(245))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(244)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(245) < ecg(244))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(244))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(245)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(244))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110101" => if(ecg(246) > ecg(245))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(246))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(245)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(246) < ecg(245))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(245))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(246)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(245))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110110" => if(ecg(247) > ecg(246))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(247))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(246)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(247) < ecg(246))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(246))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(247)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(246))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011110111" => if(ecg(248) > ecg(247))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(248))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(247)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(248) < ecg(247))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(247))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(248)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(247))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111000" => if(ecg(249) > ecg(248))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(249))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(248)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(249) < ecg(248))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(248))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(249)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(248))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111001" => if(ecg(250) > ecg(249))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(250))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(249)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(250) < ecg(249))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(249))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(250)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(249))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111010" => if(ecg(251) > ecg(250))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(251))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(250)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(251) < ecg(250))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(250))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(251)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(250))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111011" => if(ecg(252) > ecg(251))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(252))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(251)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(252) < ecg(251))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(251))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(252)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(251))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111100" => if(ecg(253) > ecg(252))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(253))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(252)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(253) < ecg(252))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(252))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(253)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(252))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111101" => if(ecg(254) > ecg(253))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(254))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(253)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(254) < ecg(253))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(253))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(254)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(253))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111110" => if(ecg(255) > ecg(254))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(255))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(254)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(255) < ecg(254))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(254))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(255)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(254))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0011111111" => if(ecg(256) > ecg(255))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(256))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(255)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(256) < ecg(255))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(255))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(256)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(255))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000000" => if(ecg(257) > ecg(256))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(257))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(256)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(257) < ecg(256))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(256))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(257)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(256))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000001" => if(ecg(258) > ecg(257))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(258))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(257)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(258) < ecg(257))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(257))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(258)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(257))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000010" => if(ecg(259) > ecg(258))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(259))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(258)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(259) < ecg(258))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(258))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(259)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(258))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000011" => if(ecg(260) > ecg(259))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(260))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(259)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(260) < ecg(259))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(259))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(260)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(259))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000100" => if(ecg(261) > ecg(260))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(261))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(260)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(261) < ecg(260))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(260))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(261)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(260))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000101" => if(ecg(262) > ecg(261))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(262))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(261)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(262) < ecg(261))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(261))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(262)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(261))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000110" => if(ecg(263) > ecg(262))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(263))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(262)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(263) < ecg(262))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(262))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(263)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(262))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100000111" => if(ecg(264) > ecg(263))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(264))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(263)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(264) < ecg(263))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(263))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(264)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(263))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001000" => if(ecg(265) > ecg(264))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(265))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(264)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(265) < ecg(264))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(264))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(265)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(264))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001001" => if(ecg(266) > ecg(265))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(266))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(265)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(266) < ecg(265))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(265))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(266)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(265))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001010" => if(ecg(267) > ecg(266))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(267))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(266)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(267) < ecg(266))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(266))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(267)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(266))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001011" => if(ecg(268) > ecg(267))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(268))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(267)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(268) < ecg(267))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(267))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(268)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(267))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001100" => if(ecg(269) > ecg(268))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(269))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(268)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(269) < ecg(268))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(268))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(269)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(268))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001101" => if(ecg(270) > ecg(269))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(270))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(269)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(270) < ecg(269))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(269))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(270)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(269))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001110" => if(ecg(271) > ecg(270))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(271))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(270)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(271) < ecg(270))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(270))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(271)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(270))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100001111" => if(ecg(272) > ecg(271))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(272))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(271)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(272) < ecg(271))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(271))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(272)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(271))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010000" => if(ecg(273) > ecg(272))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(273))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(272)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(273) < ecg(272))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(272))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(273)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(272))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010001" => if(ecg(274) > ecg(273))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(274))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(273)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(274) < ecg(273))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(273))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(274)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(273))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010010" => if(ecg(275) > ecg(274))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(275))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(274)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(275) < ecg(274))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(274))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(275)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(274))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010011" => if(ecg(276) > ecg(275))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(276))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(275)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(276) < ecg(275))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(275))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(276)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(275))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010100" => if(ecg(277) > ecg(276))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(277))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(276)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(277) < ecg(276))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(276))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(277)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(276))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010101" => if(ecg(278) > ecg(277))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(278))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(277)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(278) < ecg(277))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(277))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(278)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(277))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010110" => if(ecg(279) > ecg(278))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(279))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(278)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(279) < ecg(278))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(278))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(279)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(278))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100010111" => if(ecg(280) > ecg(279))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(280))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(279)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(280) < ecg(279))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(279))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(280)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(279))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011000" => if(ecg(281) > ecg(280))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(281))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(280)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(281) < ecg(280))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(280))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(281)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(280))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011001" => if(ecg(282) > ecg(281))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(282))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(281)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(282) < ecg(281))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(281))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(282)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(281))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011010" => if(ecg(283) > ecg(282))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(283))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(282)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(283) < ecg(282))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(282))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(283)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(282))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011011" => if(ecg(284) > ecg(283))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(284))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(283)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(284) < ecg(283))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(283))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(284)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(283))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011100" => if(ecg(285) > ecg(284))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(285))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(284)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(285) < ecg(284))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(284))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(285)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(284))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011101" => if(ecg(286) > ecg(285))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(286))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(285)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(286) < ecg(285))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(285))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(286)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(285))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011110" => if(ecg(287) > ecg(286))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(287))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(286)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(287) < ecg(286))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(286))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(287)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(286))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100011111" => if(ecg(288) > ecg(287))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(288))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(287)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(288) < ecg(287))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(287))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(288)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(287))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100000" => if(ecg(289) > ecg(288))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(289))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(288)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(289) < ecg(288))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(288))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(289)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(288))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100001" => if(ecg(290) > ecg(289))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(290))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(289)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(290) < ecg(289))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(289))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(290)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(289))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100010" => if(ecg(291) > ecg(290))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(291))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(290)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(291) < ecg(290))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(290))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(291)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(290))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100011" => if(ecg(292) > ecg(291))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(292))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(291)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(292) < ecg(291))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(291))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(292)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(291))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100100" => if(ecg(293) > ecg(292))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(293))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(292)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(293) < ecg(292))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(292))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(293)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(292))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100101" => if(ecg(294) > ecg(293))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(294))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(293)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(294) < ecg(293))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(293))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(294)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(293))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100110" => if(ecg(295) > ecg(294))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(295))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(294)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(295) < ecg(294))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(294))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(295)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(294))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100100111" => if(ecg(296) > ecg(295))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(296))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(295)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(296) < ecg(295))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(295))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(296)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(295))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101000" => if(ecg(297) > ecg(296))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(297))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(296)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(297) < ecg(296))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(296))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(297)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(296))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101001" => if(ecg(298) > ecg(297))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(298))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(297)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(298) < ecg(297))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(297))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(298)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(297))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101010" => if(ecg(299) > ecg(298))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(299))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(298)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(299) < ecg(298))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(298))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(299)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(298))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101011" => if(ecg(300) > ecg(299))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(300))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(299)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(300) < ecg(299))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(299))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(300)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(299))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101100" => if(ecg(301) > ecg(300))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(301))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(300)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(301) < ecg(300))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(300))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(301)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(300))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101101" => if(ecg(302) > ecg(301))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(302))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(301)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(302) < ecg(301))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(301))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(302)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(301))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101110" => if(ecg(303) > ecg(302))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(303))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(302)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(303) < ecg(302))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(302))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(303)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(302))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100101111" => if(ecg(304) > ecg(303))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(304))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(303)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(304) < ecg(303))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(303))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(304)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(303))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110000" => if(ecg(305) > ecg(304))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(305))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(304)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(305) < ecg(304))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(304))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(305)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(304))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110001" => if(ecg(306) > ecg(305))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(306))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(305)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(306) < ecg(305))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(305))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(306)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(305))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110010" => if(ecg(307) > ecg(306))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(307))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(306)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(307) < ecg(306))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(306))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(307)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(306))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110011" => if(ecg(308) > ecg(307))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(308))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(307)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(308) < ecg(307))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(307))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(308)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(307))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110100" => if(ecg(309) > ecg(308))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(309))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(308)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(309) < ecg(308))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(308))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(309)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(308))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110101" => if(ecg(310) > ecg(309))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(310))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(309)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(310) < ecg(309))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(309))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(310)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(309))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110110" => if(ecg(311) > ecg(310))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(311))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(310)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(311) < ecg(310))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(310))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(311)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(310))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100110111" => if(ecg(312) > ecg(311))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(312))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(311)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(312) < ecg(311))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(311))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(312)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(311))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111000" => if(ecg(313) > ecg(312))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(313))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(312)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(313) < ecg(312))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(312))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(313)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(312))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111001" => if(ecg(314) > ecg(313))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(314))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(313)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(314) < ecg(313))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(313))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(314)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(313))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111010" => if(ecg(315) > ecg(314))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(315))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(314)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(315) < ecg(314))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(314))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(315)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(314))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111011" => if(ecg(316) > ecg(315))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(316))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(315)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(316) < ecg(315))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(315))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(316)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(315))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111100" => if(ecg(317) > ecg(316))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(317))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(316)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(317) < ecg(316))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(316))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(317)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(316))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111101" => if(ecg(318) > ecg(317))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(318))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(317)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(318) < ecg(317))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(317))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(318)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(317))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111110" => if(ecg(319) > ecg(318))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(319))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(318)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(319) < ecg(318))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(318))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(319)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(318))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0100111111" => if(ecg(320) > ecg(319))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(320))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(319)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(320) < ecg(319))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(319))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(320)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(319))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000000" => if(ecg(321) > ecg(320))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(321))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(320)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(321) < ecg(320))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(320))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(321)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(320))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000001" => if(ecg(322) > ecg(321))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(322))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(321)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(322) < ecg(321))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(321))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(322)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(321))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000010" => if(ecg(323) > ecg(322))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(323))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(322)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(323) < ecg(322))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(322))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(323)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(322))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000011" => if(ecg(324) > ecg(323))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(324))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(323)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(324) < ecg(323))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(323))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(324)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(323))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000100" => if(ecg(325) > ecg(324))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(325))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(324)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(325) < ecg(324))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(324))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(325)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(324))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000101" => if(ecg(326) > ecg(325))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(326))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(325)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(326) < ecg(325))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(325))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(326)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(325))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000110" => if(ecg(327) > ecg(326))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(327))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(326)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(327) < ecg(326))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(326))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(327)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(326))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101000111" => if(ecg(328) > ecg(327))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(328))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(327)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(328) < ecg(327))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(327))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(328)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(327))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001000" => if(ecg(329) > ecg(328))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(329))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(328)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(329) < ecg(328))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(328))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(329)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(328))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001001" => if(ecg(330) > ecg(329))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(330))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(329)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(330) < ecg(329))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(329))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(330)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(329))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001010" => if(ecg(331) > ecg(330))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(331))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(330)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(331) < ecg(330))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(330))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(331)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(330))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001011" => if(ecg(332) > ecg(331))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(332))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(331)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(332) < ecg(331))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(331))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(332)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(331))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001100" => if(ecg(333) > ecg(332))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(333))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(332)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(333) < ecg(332))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(332))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(333)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(332))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001101" => if(ecg(334) > ecg(333))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(334))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(333)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(334) < ecg(333))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(333))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(334)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(333))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001110" => if(ecg(335) > ecg(334))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(335))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(334)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(335) < ecg(334))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(334))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(335)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(334))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101001111" => if(ecg(336) > ecg(335))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(336))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(335)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(336) < ecg(335))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(335))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(336)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(335))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010000" => if(ecg(337) > ecg(336))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(337))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(336)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(337) < ecg(336))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(336))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(337)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(336))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010001" => if(ecg(338) > ecg(337))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(338))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(337)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(338) < ecg(337))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(337))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(338)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(337))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010010" => if(ecg(339) > ecg(338))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(339))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(338)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(339) < ecg(338))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(338))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(339)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(338))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010011" => if(ecg(340) > ecg(339))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(340))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(339)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(340) < ecg(339))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(339))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(340)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(339))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010100" => if(ecg(341) > ecg(340))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(341))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(340)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(341) < ecg(340))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(340))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(341)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(340))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010101" => if(ecg(342) > ecg(341))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(342))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(341)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(342) < ecg(341))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(341))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(342)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(341))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010110" => if(ecg(343) > ecg(342))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(343))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(342)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(343) < ecg(342))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(342))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(343)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(342))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101010111" => if(ecg(344) > ecg(343))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(344))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(343)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(344) < ecg(343))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(343))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(344)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(343))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011000" => if(ecg(345) > ecg(344))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(345))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(344)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(345) < ecg(344))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(344))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(345)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(344))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011001" => if(ecg(346) > ecg(345))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(346))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(345)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(346) < ecg(345))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(345))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(346)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(345))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011010" => if(ecg(347) > ecg(346))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(347))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(346)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(347) < ecg(346))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(346))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(347)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(346))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011011" => if(ecg(348) > ecg(347))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(348))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(347)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(348) < ecg(347))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(347))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(348)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(347))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011100" => if(ecg(349) > ecg(348))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(349))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(348)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(349) < ecg(348))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(348))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(349)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(348))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011101" => if(ecg(350) > ecg(349))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(350))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(349)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(350) < ecg(349))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(349))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(350)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(349))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011110" => if(ecg(351) > ecg(350))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(351))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(350)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(351) < ecg(350))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(350))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(351)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(350))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101011111" => if(ecg(352) > ecg(351))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(352))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(351)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(352) < ecg(351))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(351))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(352)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(351))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100000" => if(ecg(353) > ecg(352))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(353))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(352)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(353) < ecg(352))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(352))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(353)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(352))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100001" => if(ecg(354) > ecg(353))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(354))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(353)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(354) < ecg(353))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(353))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(354)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(353))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100010" => if(ecg(355) > ecg(354))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(355))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(354)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(355) < ecg(354))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(354))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(355)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(354))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100011" => if(ecg(356) > ecg(355))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(356))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(355)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(356) < ecg(355))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(355))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(356)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(355))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100100" => if(ecg(357) > ecg(356))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(357))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(356)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(357) < ecg(356))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(356))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(357)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(356))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100101" => if(ecg(358) > ecg(357))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(358))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(357)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(358) < ecg(357))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(357))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(358)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(357))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100110" => if(ecg(359) > ecg(358))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(359))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(358)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(359) < ecg(358))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(358))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(359)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(358))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101100111" => if(ecg(360) > ecg(359))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(360))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(359)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(360) < ecg(359))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(359))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(360)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(359))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101000" => if(ecg(361) > ecg(360))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(361))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(360)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(361) < ecg(360))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(360))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(361)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(360))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101001" => if(ecg(362) > ecg(361))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(362))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(361)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(362) < ecg(361))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(361))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(362)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(361))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101010" => if(ecg(363) > ecg(362))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(363))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(362)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(363) < ecg(362))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(362))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(363)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(362))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101011" => if(ecg(364) > ecg(363))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(364))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(363)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(364) < ecg(363))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(363))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(364)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(363))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101100" => if(ecg(365) > ecg(364))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(365))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(364)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(365) < ecg(364))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(364))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(365)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(364))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101101" => if(ecg(366) > ecg(365))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(366))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(365)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(366) < ecg(365))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(365))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(366)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(365))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101110" => if(ecg(367) > ecg(366))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(367))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(366)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(367) < ecg(366))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(366))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(367)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(366))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101101111" => if(ecg(368) > ecg(367))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(368))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(367)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(368) < ecg(367))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(367))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(368)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(367))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110000" => if(ecg(369) > ecg(368))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(369))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(368)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(369) < ecg(368))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(368))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(369)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(368))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110001" => if(ecg(370) > ecg(369))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(370))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(369)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(370) < ecg(369))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(369))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(370)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(369))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110010" => if(ecg(371) > ecg(370))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(371))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(370)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(371) < ecg(370))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(370))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(371)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(370))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110011" => if(ecg(372) > ecg(371))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(372))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(371)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(372) < ecg(371))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(371))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(372)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(371))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110100" => if(ecg(373) > ecg(372))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(373))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(372)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(373) < ecg(372))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(372))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(373)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(372))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110101" => if(ecg(374) > ecg(373))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(374))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(373)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(374) < ecg(373))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(373))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(374)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(373))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110110" => if(ecg(375) > ecg(374))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(375))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(374)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(375) < ecg(374))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(374))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(375)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(374))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101110111" => if(ecg(376) > ecg(375))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(376))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(375)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(376) < ecg(375))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(375))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(376)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(375))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111000" => if(ecg(377) > ecg(376))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(377))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(376)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(377) < ecg(376))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(376))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(377)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(376))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111001" => if(ecg(378) > ecg(377))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(378))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(377)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(378) < ecg(377))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(377))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(378)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(377))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111010" => if(ecg(379) > ecg(378))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(379))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(378)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(379) < ecg(378))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(378))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(379)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(378))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111011" => if(ecg(380) > ecg(379))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(380))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(379)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(380) < ecg(379))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(379))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(380)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(379))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111100" => if(ecg(381) > ecg(380))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(381))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(380)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(381) < ecg(380))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(380))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(381)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(380))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111101" => if(ecg(382) > ecg(381))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(382))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(381)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(382) < ecg(381))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(381))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(382)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(381))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111110" => if(ecg(383) > ecg(382))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(383))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(382)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(383) < ecg(382))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(382))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(383)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(382))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0101111111" => if(ecg(384) > ecg(383))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(384))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(383)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(384) < ecg(383))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(383))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(384)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(383))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000000" => if(ecg(385) > ecg(384))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(385))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(384)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(385) < ecg(384))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(384))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(385)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(384))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000001" => if(ecg(386) > ecg(385))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(386))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(385)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(386) < ecg(385))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(385))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(386)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(385))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000010" => if(ecg(387) > ecg(386))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(387))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(386)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(387) < ecg(386))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(386))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(387)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(386))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000011" => if(ecg(388) > ecg(387))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(388))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(387)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(388) < ecg(387))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(387))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(388)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(387))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000100" => if(ecg(389) > ecg(388))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(389))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(388)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(389) < ecg(388))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(388))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(389)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(388))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000101" => if(ecg(390) > ecg(389))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(390))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(389)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(390) < ecg(389))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(389))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(390)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(389))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000110" => if(ecg(391) > ecg(390))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(391))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(390)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(391) < ecg(390))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(390))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(391)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(390))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110000111" => if(ecg(392) > ecg(391))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(392))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(391)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(392) < ecg(391))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(391))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(392)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(391))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001000" => if(ecg(393) > ecg(392))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(393))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(392)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(393) < ecg(392))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(392))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(393)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(392))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001001" => if(ecg(394) > ecg(393))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(394))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(393)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(394) < ecg(393))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(393))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(394)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(393))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001010" => if(ecg(395) > ecg(394))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(395))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(394)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(395) < ecg(394))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(394))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(395)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(394))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001011" => if(ecg(396) > ecg(395))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(396))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(395)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(396) < ecg(395))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(395))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(396)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(395))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001100" => if(ecg(397) > ecg(396))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(397))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(396)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(397) < ecg(396))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(396))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(397)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(396))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001101" => if(ecg(398) > ecg(397))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(398))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(397)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(398) < ecg(397))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(397))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(398)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(397))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001110" => if(ecg(399) > ecg(398))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(399))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(398)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(399) < ecg(398))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(398))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(399)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(398))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110001111" => if(ecg(400) > ecg(399))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(400))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(399)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(400) < ecg(399))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(399))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(400)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(399))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010000" => if(ecg(401) > ecg(400))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(401))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(400)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(401) < ecg(400))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(400))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(401)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(400))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010001" => if(ecg(402) > ecg(401))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(402))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(401)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(402) < ecg(401))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(401))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(402)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(401))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010010" => if(ecg(403) > ecg(402))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(403))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(402)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(403) < ecg(402))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(402))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(403)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(402))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010011" => if(ecg(404) > ecg(403))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(404))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(403)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(404) < ecg(403))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(403))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(404)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(403))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010100" => if(ecg(405) > ecg(404))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(405))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(404)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(405) < ecg(404))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(404))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(405)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(404))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010101" => if(ecg(406) > ecg(405))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(406))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(405)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(406) < ecg(405))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(405))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(406)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(405))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010110" => if(ecg(407) > ecg(406))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(407))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(406)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(407) < ecg(406))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(406))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(407)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(406))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110010111" => if(ecg(408) > ecg(407))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(408))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(407)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(408) < ecg(407))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(407))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(408)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(407))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011000" => if(ecg(409) > ecg(408))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(409))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(408)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(409) < ecg(408))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(408))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(409)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(408))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011001" => if(ecg(410) > ecg(409))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(410))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(409)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(410) < ecg(409))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(409))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(410)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(409))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011010" => if(ecg(411) > ecg(410))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(411))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(410)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(411) < ecg(410))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(410))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(411)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(410))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011011" => if(ecg(412) > ecg(411))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(412))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(411)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(412) < ecg(411))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(411))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(412)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(411))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011100" => if(ecg(413) > ecg(412))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(413))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(412)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(413) < ecg(412))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(412))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(413)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(412))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011101" => if(ecg(414) > ecg(413))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(414))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(413)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(414) < ecg(413))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(413))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(414)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(413))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011110" => if(ecg(415) > ecg(414))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(415))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(414)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(415) < ecg(414))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(414))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(415)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(414))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110011111" => if(ecg(416) > ecg(415))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(416))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(415)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(416) < ecg(415))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(415))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(416)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(415))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100000" => if(ecg(417) > ecg(416))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(417))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(416)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(417) < ecg(416))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(416))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(417)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(416))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100001" => if(ecg(418) > ecg(417))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(418))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(417)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(418) < ecg(417))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(417))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(418)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(417))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100010" => if(ecg(419) > ecg(418))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(419))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(418)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(419) < ecg(418))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(418))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(419)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(418))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100011" => if(ecg(420) > ecg(419))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(420))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(419)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(420) < ecg(419))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(419))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(420)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(419))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100100" => if(ecg(421) > ecg(420))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(421))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(420)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(421) < ecg(420))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(420))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(421)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(420))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100101" => if(ecg(422) > ecg(421))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(422))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(421)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(422) < ecg(421))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(421))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(422)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(421))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100110" => if(ecg(423) > ecg(422))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(423))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(422)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(423) < ecg(422))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(422))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(423)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(422))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110100111" => if(ecg(424) > ecg(423))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(424))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(423)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(424) < ecg(423))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(423))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(424)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(423))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101000" => if(ecg(425) > ecg(424))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(425))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(424)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(425) < ecg(424))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(424))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(425)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(424))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101001" => if(ecg(426) > ecg(425))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(426))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(425)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(426) < ecg(425))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(425))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(426)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(425))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101010" => if(ecg(427) > ecg(426))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(427))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(426)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(427) < ecg(426))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(426))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(427)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(426))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101011" => if(ecg(428) > ecg(427))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(428))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(427)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(428) < ecg(427))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(427))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(428)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(427))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101100" => if(ecg(429) > ecg(428))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(429))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(428)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(429) < ecg(428))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(428))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(429)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(428))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101101" => if(ecg(430) > ecg(429))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(430))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(429)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(430) < ecg(429))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(429))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(430)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(429))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101110" => if(ecg(431) > ecg(430))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(431))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(430)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(431) < ecg(430))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(430))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(431)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(430))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110101111" => if(ecg(432) > ecg(431))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(432))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(431)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(432) < ecg(431))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(431))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(432)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(431))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110000" => if(ecg(433) > ecg(432))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(433))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(432)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(433) < ecg(432))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(432))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(433)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(432))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110001" => if(ecg(434) > ecg(433))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(434))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(433)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(434) < ecg(433))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(433))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(434)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(433))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110010" => if(ecg(435) > ecg(434))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(435))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(434)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(435) < ecg(434))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(434))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(435)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(434))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110011" => if(ecg(436) > ecg(435))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(436))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(435)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(436) < ecg(435))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(435))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(436)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(435))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110100" => if(ecg(437) > ecg(436))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(437))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(436)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(437) < ecg(436))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(436))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(437)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(436))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110101" => if(ecg(438) > ecg(437))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(438))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(437)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(438) < ecg(437))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(437))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(438)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(437))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110110" => if(ecg(439) > ecg(438))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(439))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(438)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(439) < ecg(438))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(438))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(439)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(438))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110110111" => if(ecg(440) > ecg(439))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(440))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(439)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(440) < ecg(439))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(439))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(440)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(439))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111000" => if(ecg(441) > ecg(440))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(441))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(440)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(441) < ecg(440))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(440))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(441)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(440))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111001" => if(ecg(442) > ecg(441))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(442))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(441)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(442) < ecg(441))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(441))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(442)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(441))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111010" => if(ecg(443) > ecg(442))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(443))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(442)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(443) < ecg(442))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(442))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(443)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(442))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111011" => if(ecg(444) > ecg(443))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(444))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(443)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(444) < ecg(443))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(443))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(444)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(443))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111100" => if(ecg(445) > ecg(444))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(445))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(444)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(445) < ecg(444))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(444))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(445)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(444))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111101" => if(ecg(446) > ecg(445))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(446))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(445)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(446) < ecg(445))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(445))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(446)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(445))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111110" => if(ecg(447) > ecg(446))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(447))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(446)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(447) < ecg(446))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(446))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(447)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(446))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0110111111" => if(ecg(448) > ecg(447))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(448))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(447)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(448) < ecg(447))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(447))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(448)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(447))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000000" => if(ecg(449) > ecg(448))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(449))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(448)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(449) < ecg(448))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(448))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(449)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(448))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000001" => if(ecg(450) > ecg(449))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(450))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(449)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(450) < ecg(449))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(449))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(450)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(449))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000010" => if(ecg(451) > ecg(450))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(451))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(450)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(451) < ecg(450))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(450))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(451)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(450))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000011" => if(ecg(452) > ecg(451))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(452))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(451)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(452) < ecg(451))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(451))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(452)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(451))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000100" => if(ecg(453) > ecg(452))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(453))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(452)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(453) < ecg(452))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(452))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(453)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(452))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000101" => if(ecg(454) > ecg(453))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(454))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(453)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(454) < ecg(453))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(453))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(454)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(453))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000110" => if(ecg(455) > ecg(454))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(455))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(454)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(455) < ecg(454))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(454))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(455)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(454))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111000111" => if(ecg(456) > ecg(455))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(456))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(455)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(456) < ecg(455))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(455))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(456)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(455))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001000" => if(ecg(457) > ecg(456))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(457))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(456)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(457) < ecg(456))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(456))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(457)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(456))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001001" => if(ecg(458) > ecg(457))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(458))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(457)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(458) < ecg(457))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(457))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(458)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(457))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001010" => if(ecg(459) > ecg(458))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(459))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(458)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(459) < ecg(458))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(458))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(459)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(458))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001011" => if(ecg(460) > ecg(459))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(460))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(459)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(460) < ecg(459))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(459))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(460)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(459))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001100" => if(ecg(461) > ecg(460))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(461))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(460)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(461) < ecg(460))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(460))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(461)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(460))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001101" => if(ecg(462) > ecg(461))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(462))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(461)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(462) < ecg(461))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(461))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(462)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(461))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001110" => if(ecg(463) > ecg(462))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(463))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(462)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(463) < ecg(462))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(462))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(463)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(462))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111001111" => if(ecg(464) > ecg(463))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(464))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(463)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(464) < ecg(463))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(463))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(464)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(463))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010000" => if(ecg(465) > ecg(464))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(465))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(464)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(465) < ecg(464))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(464))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(465)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(464))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010001" => if(ecg(466) > ecg(465))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(466))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(465)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(466) < ecg(465))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(465))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(466)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(465))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010010" => if(ecg(467) > ecg(466))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(467))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(466)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(467) < ecg(466))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(466))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(467)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(466))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010011" => if(ecg(468) > ecg(467))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(468))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(467)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(468) < ecg(467))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(467))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(468)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(467))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010100" => if(ecg(469) > ecg(468))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(469))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(468)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(469) < ecg(468))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(468))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(469)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(468))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010101" => if(ecg(470) > ecg(469))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(470))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(469)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(470) < ecg(469))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(469))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(470)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(469))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010110" => if(ecg(471) > ecg(470))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(471))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(470)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(471) < ecg(470))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(470))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(471)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(470))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111010111" => if(ecg(472) > ecg(471))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(472))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(471)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(472) < ecg(471))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(471))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(472)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(471))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011000" => if(ecg(473) > ecg(472))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(473))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(472)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(473) < ecg(472))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(472))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(473)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(472))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011001" => if(ecg(474) > ecg(473))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(474))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(473)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(474) < ecg(473))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(473))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(474)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(473))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011010" => if(ecg(475) > ecg(474))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(475))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(474)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(475) < ecg(474))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(474))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(475)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(474))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011011" => if(ecg(476) > ecg(475))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(476))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(475)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(476) < ecg(475))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(475))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(476)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(475))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011100" => if(ecg(477) > ecg(476))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(477))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(476)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(477) < ecg(476))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(476))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(477)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(476))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011101" => if(ecg(478) > ecg(477))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(478))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(477)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(478) < ecg(477))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(477))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(478)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(477))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011110" => if(ecg(479) > ecg(478))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(479))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(478)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(479) < ecg(478))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(478))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(479)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(478))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111011111" => if(ecg(480) > ecg(479))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(480))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(479)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(480) < ecg(479))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(479))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(480)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(479))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100000" => if(ecg(481) > ecg(480))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(481))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(480)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(481) < ecg(480))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(480))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(481)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(480))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100001" => if(ecg(482) > ecg(481))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(482))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(481)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(482) < ecg(481))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(481))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(482)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(481))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100010" => if(ecg(483) > ecg(482))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(483))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(482)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(483) < ecg(482))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(482))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(483)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(482))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100011" => if(ecg(484) > ecg(483))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(484))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(483)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(484) < ecg(483))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(483))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(484)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(483))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100100" => if(ecg(485) > ecg(484))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(485))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(484)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(485) < ecg(484))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(484))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(485)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(484))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100101" => if(ecg(486) > ecg(485))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(486))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(485)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(486) < ecg(485))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(485))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(486)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(485))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100110" => if(ecg(487) > ecg(486))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(487))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(486)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(487) < ecg(486))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(486))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(487)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(486))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111100111" => if(ecg(488) > ecg(487))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(488))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(487)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(488) < ecg(487))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(487))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(488)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(487))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101000" => if(ecg(489) > ecg(488))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(489))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(488)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(489) < ecg(488))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(488))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(489)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(488))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101001" => if(ecg(490) > ecg(489))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(490))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(489)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(490) < ecg(489))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(489))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(490)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(489))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101010" => if(ecg(491) > ecg(490))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(491))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(490)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(491) < ecg(490))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(490))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(491)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(490))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101011" => if(ecg(492) > ecg(491))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(492))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(491)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(492) < ecg(491))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(491))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(492)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(491))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101100" => if(ecg(493) > ecg(492))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(493))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(492)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(493) < ecg(492))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(492))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(493)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(492))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101101" => if(ecg(494) > ecg(493))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(494))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(493)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(494) < ecg(493))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(493))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(494)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(493))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101110" => if(ecg(495) > ecg(494))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(495))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(494)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(495) < ecg(494))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(494))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(495)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(494))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111101111" => if(ecg(496) > ecg(495))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(496))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(495)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(496) < ecg(495))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(495))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(496)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(495))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110000" => if(ecg(497) > ecg(496))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(497))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(496)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(497) < ecg(496))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(496))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(497)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(496))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110001" => if(ecg(498) > ecg(497))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(498))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(497)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(498) < ecg(497))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(497))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(498)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(497))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110010" => if(ecg(499) > ecg(498))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(499))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(498)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(499) < ecg(498))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(498))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(499)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(498))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110011" => if(ecg(500) > ecg(499))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(500))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(499)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(500) < ecg(499))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(499))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(500)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(499))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110100" => if(ecg(501) > ecg(500))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(501))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(500)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(501) < ecg(500))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(500))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(501)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(500))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110101" => if(ecg(502) > ecg(501))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(502))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(501)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(502) < ecg(501))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(501))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(502)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(501))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110110" => if(ecg(503) > ecg(502))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(503))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(502)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(503) < ecg(502))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(502))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(503)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(502))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111110111" => if(ecg(504) > ecg(503))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(504))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(503)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(504) < ecg(503))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(503))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(504)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(503))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111000" => if(ecg(505) > ecg(504))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(505))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(504)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(505) < ecg(504))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(504))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(505)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(504))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111001" => if(ecg(506) > ecg(505))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(506))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(505)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(506) < ecg(505))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(505))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(506)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(505))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111010" => if(ecg(507) > ecg(506))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(507))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(506)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(507) < ecg(506))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(506))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(507)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(506))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111011" => if(ecg(508) > ecg(507))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(508))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(507)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(508) < ecg(507))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(507))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(508)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(507))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111100" => if(ecg(509) > ecg(508))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(509))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(508)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(509) < ecg(508))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(508))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(509)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(508))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111101" => if(ecg(510) > ecg(509))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(510))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(509)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(510) < ecg(509))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(509))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(510)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(509))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111110" => if(ecg(511) > ecg(510))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(511))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(510)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(511) < ecg(510))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(510))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(511)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(510))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "0111111111" => if(ecg(512) > ecg(511))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(512))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(511)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(512) < ecg(511))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(511))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(512)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(511))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000000" => if(ecg(513) > ecg(512))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(513))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(512)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(513) < ecg(512))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(512))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(513)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(512))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000001" => if(ecg(514) > ecg(513))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(514))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(513)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(514) < ecg(513))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(513))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(514)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(513))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000010" => if(ecg(515) > ecg(514))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(515))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(514)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(515) < ecg(514))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(514))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(515)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(514))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000011" => if(ecg(516) > ecg(515))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(516))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(515)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(516) < ecg(515))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(515))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(516)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(515))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000100" => if(ecg(517) > ecg(516))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(517))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(516)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(517) < ecg(516))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(516))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(517)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(516))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000101" => if(ecg(518) > ecg(517))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(518))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(517)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(518) < ecg(517))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(517))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(518)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(517))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000110" => if(ecg(519) > ecg(518))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(519))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(518)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(519) < ecg(518))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(518))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(519)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(518))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000000111" => if(ecg(520) > ecg(519))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(520))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(519)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(520) < ecg(519))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(519))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(520)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(519))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001000" => if(ecg(521) > ecg(520))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(521))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(520)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(521) < ecg(520))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(520))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(521)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(520))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001001" => if(ecg(522) > ecg(521))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(522))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(521)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(522) < ecg(521))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(521))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(522)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(521))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001010" => if(ecg(523) > ecg(522))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(523))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(522)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(523) < ecg(522))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(522))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(523)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(522))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001011" => if(ecg(524) > ecg(523))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(524))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(523)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(524) < ecg(523))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(523))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(524)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(523))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001100" => if(ecg(525) > ecg(524))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(525))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(524)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(525) < ecg(524))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(524))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(525)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(524))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001101" => if(ecg(526) > ecg(525))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(526))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(525)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(526) < ecg(525))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(525))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(526)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(525))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001110" => if(ecg(527) > ecg(526))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(527))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(526)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(527) < ecg(526))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(526))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(527)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(526))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000001111" => if(ecg(528) > ecg(527))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(528))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(527)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(528) < ecg(527))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(527))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(528)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(527))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010000" => if(ecg(529) > ecg(528))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(529))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(528)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(529) < ecg(528))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(528))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(529)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(528))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010001" => if(ecg(530) > ecg(529))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(530))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(529)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(530) < ecg(529))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(529))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(530)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(529))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010010" => if(ecg(531) > ecg(530))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(531))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(530)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(531) < ecg(530))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(530))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(531)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(530))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010011" => if(ecg(532) > ecg(531))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(532))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(531)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(532) < ecg(531))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(531))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(532)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(531))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010100" => if(ecg(533) > ecg(532))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(533))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(532)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(533) < ecg(532))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(532))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(533)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(532))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010101" => if(ecg(534) > ecg(533))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(534))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(533)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(534) < ecg(533))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(533))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(534)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(533))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010110" => if(ecg(535) > ecg(534))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(535))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(534)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(535) < ecg(534))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(534))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(535)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(534))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000010111" => if(ecg(536) > ecg(535))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(536))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(535)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(536) < ecg(535))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(535))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(536)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(535))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011000" => if(ecg(537) > ecg(536))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(537))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(536)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(537) < ecg(536))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(536))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(537)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(536))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011001" => if(ecg(538) > ecg(537))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(538))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(537)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(538) < ecg(537))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(537))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(538)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(537))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011010" => if(ecg(539) > ecg(538))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(539))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(538)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(539) < ecg(538))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(538))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(539)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(538))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011011" => if(ecg(540) > ecg(539))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(540))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(539)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(540) < ecg(539))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(539))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(540)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(539))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011100" => if(ecg(541) > ecg(540))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(541))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(540)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(541) < ecg(540))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(540))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(541)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(540))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011101" => if(ecg(542) > ecg(541))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(542))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(541)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(542) < ecg(541))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(541))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(542)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(541))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011110" => if(ecg(543) > ecg(542))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(543))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(542)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(543) < ecg(542))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(542))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(543)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(542))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000011111" => if(ecg(544) > ecg(543))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(544))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(543)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(544) < ecg(543))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(543))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(544)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(543))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100000" => if(ecg(545) > ecg(544))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(545))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(544)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(545) < ecg(544))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(544))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(545)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(544))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100001" => if(ecg(546) > ecg(545))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(546))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(545)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(546) < ecg(545))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(545))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(546)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(545))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100010" => if(ecg(547) > ecg(546))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(547))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(546)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(547) < ecg(546))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(546))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(547)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(546))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100011" => if(ecg(548) > ecg(547))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(548))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(547)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(548) < ecg(547))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(547))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(548)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(547))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100100" => if(ecg(549) > ecg(548))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(549))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(548)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(549) < ecg(548))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(548))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(549)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(548))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100101" => if(ecg(550) > ecg(549))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(550))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(549)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(550) < ecg(549))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(549))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(550)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(549))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100110" => if(ecg(551) > ecg(550))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(551))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(550)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(551) < ecg(550))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(550))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(551)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(550))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000100111" => if(ecg(552) > ecg(551))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(552))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(551)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(552) < ecg(551))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(551))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(552)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(551))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101000" => if(ecg(553) > ecg(552))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(553))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(552)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(553) < ecg(552))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(552))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(553)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(552))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101001" => if(ecg(554) > ecg(553))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(554))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(553)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(554) < ecg(553))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(553))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(554)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(553))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101010" => if(ecg(555) > ecg(554))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(555))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(554)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(555) < ecg(554))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(554))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(555)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(554))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101011" => if(ecg(556) > ecg(555))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(556))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(555)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(556) < ecg(555))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(555))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(556)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(555))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101100" => if(ecg(557) > ecg(556))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(557))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(556)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(557) < ecg(556))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(556))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(557)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(556))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101101" => if(ecg(558) > ecg(557))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(558))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(557)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(558) < ecg(557))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(557))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(558)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(557))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101110" => if(ecg(559) > ecg(558))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(559))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(558)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(559) < ecg(558))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(558))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(559)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(558))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000101111" => if(ecg(560) > ecg(559))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(560))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(559)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(560) < ecg(559))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(559))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(560)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(559))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110000" => if(ecg(561) > ecg(560))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(561))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(560)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(561) < ecg(560))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(560))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(561)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(560))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110001" => if(ecg(562) > ecg(561))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(562))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(561)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(562) < ecg(561))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(561))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(562)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(561))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110010" => if(ecg(563) > ecg(562))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(563))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(562)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(563) < ecg(562))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(562))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(563)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(562))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110011" => if(ecg(564) > ecg(563))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(564))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(563)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(564) < ecg(563))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(563))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(564)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(563))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110100" => if(ecg(565) > ecg(564))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(565))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(564)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(565) < ecg(564))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(564))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(565)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(564))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110101" => if(ecg(566) > ecg(565))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(566))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(565)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(566) < ecg(565))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(565))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(566)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(565))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110110" => if(ecg(567) > ecg(566))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(567))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(566)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(567) < ecg(566))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(566))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(567)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(566))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000110111" => if(ecg(568) > ecg(567))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(568))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(567)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(568) < ecg(567))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(567))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(568)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(567))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111000" => if(ecg(569) > ecg(568))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(569))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(568)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(569) < ecg(568))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(568))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(569)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(568))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111001" => if(ecg(570) > ecg(569))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(570))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(569)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(570) < ecg(569))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(569))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(570)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(569))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111010" => if(ecg(571) > ecg(570))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(571))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(570)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(571) < ecg(570))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(570))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(571)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(570))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111011" => if(ecg(572) > ecg(571))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(572))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(571)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(572) < ecg(571))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(571))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(572)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(571))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111100" => if(ecg(573) > ecg(572))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(573))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(572)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(573) < ecg(572))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(572))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(573)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(572))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111101" => if(ecg(574) > ecg(573))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(574))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(573)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(574) < ecg(573))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(573))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(574)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(573))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111110" => if(ecg(575) > ecg(574))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(575))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(574)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(575) < ecg(574))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(574))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(575)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(574))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1000111111" => if(ecg(576) > ecg(575))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(576))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(575)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(576) < ecg(575))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(575))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(576)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(575))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000000" => if(ecg(577) > ecg(576))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(577))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(576)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(577) < ecg(576))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(576))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(577)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(576))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000001" => if(ecg(578) > ecg(577))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(578))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(577)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(578) < ecg(577))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(577))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(578)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(577))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000010" => if(ecg(579) > ecg(578))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(579))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(578)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(579) < ecg(578))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(578))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(579)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(578))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000011" => if(ecg(580) > ecg(579))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(580))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(579)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(580) < ecg(579))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(579))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(580)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(579))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000100" => if(ecg(581) > ecg(580))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(581))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(580)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(581) < ecg(580))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(580))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(581)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(580))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000101" => if(ecg(582) > ecg(581))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(582))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(581)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(582) < ecg(581))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(581))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(582)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(581))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000110" => if(ecg(583) > ecg(582))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(583))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(582)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(583) < ecg(582))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(582))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(583)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(582))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001000111" => if(ecg(584) > ecg(583))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(584))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(583)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(584) < ecg(583))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(583))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(584)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(583))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001000" => if(ecg(585) > ecg(584))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(585))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(584)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(585) < ecg(584))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(584))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(585)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(584))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001001" => if(ecg(586) > ecg(585))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(586))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(585)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(586) < ecg(585))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(585))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(586)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(585))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001010" => if(ecg(587) > ecg(586))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(587))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(586)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(587) < ecg(586))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(586))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(587)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(586))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001011" => if(ecg(588) > ecg(587))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(588))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(587)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(588) < ecg(587))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(587))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(588)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(587))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001100" => if(ecg(589) > ecg(588))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(589))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(588)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(589) < ecg(588))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(588))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(589)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(588))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001101" => if(ecg(590) > ecg(589))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(590))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(589)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(590) < ecg(589))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(589))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(590)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(589))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001110" => if(ecg(591) > ecg(590))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(591))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(590)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(591) < ecg(590))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(590))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(591)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(590))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001001111" => if(ecg(592) > ecg(591))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(592))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(591)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(592) < ecg(591))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(591))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(592)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(591))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010000" => if(ecg(593) > ecg(592))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(593))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(592)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(593) < ecg(592))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(592))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(593)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(592))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010001" => if(ecg(594) > ecg(593))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(594))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(593)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(594) < ecg(593))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(593))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(594)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(593))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010010" => if(ecg(595) > ecg(594))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(595))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(594)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(595) < ecg(594))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(594))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(595)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(594))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010011" => if(ecg(596) > ecg(595))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(596))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(595)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(596) < ecg(595))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(595))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(596)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(595))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010100" => if(ecg(597) > ecg(596))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(597))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(596)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(597) < ecg(596))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(596))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(597)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(596))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010101" => if(ecg(598) > ecg(597))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(598))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(597)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(598) < ecg(597))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(597))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(598)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(597))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010110" => if(ecg(599) > ecg(598))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(599))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(598)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(599) < ecg(598))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(598))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(599)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(598))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001010111" => if(ecg(600) > ecg(599))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(600))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(599)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(600) < ecg(599))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(599))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(600)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(599))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011000" => if(ecg(601) > ecg(600))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(601))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(600)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(601) < ecg(600))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(600))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(601)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(600))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011001" => if(ecg(602) > ecg(601))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(602))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(601)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(602) < ecg(601))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(601))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(602)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(601))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011010" => if(ecg(603) > ecg(602))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(603))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(602)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(603) < ecg(602))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(602))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(603)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(602))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011011" => if(ecg(604) > ecg(603))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(604))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(603)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(604) < ecg(603))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(603))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(604)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(603))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011100" => if(ecg(605) > ecg(604))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(605))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(604)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(605) < ecg(604))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(604))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(605)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(604))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011101" => if(ecg(606) > ecg(605))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(606))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(605)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(606) < ecg(605))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(605))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(606)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(605))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011110" => if(ecg(607) > ecg(606))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(607))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(606)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(607) < ecg(606))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(606))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(607)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(606))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001011111" => if(ecg(608) > ecg(607))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(608))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(607)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(608) < ecg(607))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(607))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(608)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(607))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100000" => if(ecg(609) > ecg(608))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(609))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(608)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(609) < ecg(608))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(608))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(609)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(608))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100001" => if(ecg(610) > ecg(609))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(610))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(609)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(610) < ecg(609))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(609))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(610)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(609))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100010" => if(ecg(611) > ecg(610))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(611))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(610)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(611) < ecg(610))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(610))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(611)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(610))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100011" => if(ecg(612) > ecg(611))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(612))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(611)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(612) < ecg(611))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(611))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(612)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(611))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100100" => if(ecg(613) > ecg(612))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(613))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(612)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(613) < ecg(612))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(612))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(613)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(612))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100101" => if(ecg(614) > ecg(613))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(614))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(613)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(614) < ecg(613))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(613))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(614)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(613))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100110" => if(ecg(615) > ecg(614))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(615))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(614)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(615) < ecg(614))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(614))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(615)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(614))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001100111" => if(ecg(616) > ecg(615))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(616))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(615)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(616) < ecg(615))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(615))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(616)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(615))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101000" => if(ecg(617) > ecg(616))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(617))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(616)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(617) < ecg(616))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(616))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(617)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(616))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101001" => if(ecg(618) > ecg(617))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(618))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(617)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(618) < ecg(617))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(617))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(618)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(617))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101010" => if(ecg(619) > ecg(618))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(619))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(618)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(619) < ecg(618))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(618))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(619)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(618))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101011" => if(ecg(620) > ecg(619))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(620))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(619)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(620) < ecg(619))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(619))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(620)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(619))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101100" => if(ecg(621) > ecg(620))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(621))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(620)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(621) < ecg(620))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(620))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(621)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(620))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101101" => if(ecg(622) > ecg(621))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(622))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(621)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(622) < ecg(621))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(621))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(622)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(621))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101110" => if(ecg(623) > ecg(622))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(623))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(622)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(623) < ecg(622))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(622))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(623)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(622))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001101111" => if(ecg(624) > ecg(623))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(624))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(623)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(624) < ecg(623))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(623))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(624)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(623))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110000" => if(ecg(625) > ecg(624))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(625))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(624)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(625) < ecg(624))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(624))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(625)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(624))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110001" => if(ecg(626) > ecg(625))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(626))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(625)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(626) < ecg(625))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(625))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(626)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(625))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110010" => if(ecg(627) > ecg(626))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(627))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(626)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(627) < ecg(626))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(626))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(627)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(626))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110011" => if(ecg(628) > ecg(627))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(628))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(627)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(628) < ecg(627))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(627))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(628)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(627))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110100" => if(ecg(629) > ecg(628))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(629))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(628)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(629) < ecg(628))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(628))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(629)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(628))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110101" => if(ecg(630) > ecg(629))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(630))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(629)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(630) < ecg(629))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(629))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(630)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(629))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110110" => if(ecg(631) > ecg(630))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(631))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(630)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(631) < ecg(630))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(630))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(631)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(630))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001110111" => if(ecg(632) > ecg(631))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(632))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(631)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(632) < ecg(631))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(631))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(632)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(631))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111000" => if(ecg(633) > ecg(632))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(633))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(632)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(633) < ecg(632))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(632))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(633)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(632))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111001" => if(ecg(634) > ecg(633))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(634))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(633)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(634) < ecg(633))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(633))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(634)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(633))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111010" => if(ecg(635) > ecg(634))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(635))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(634)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(635) < ecg(634))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(634))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(635)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(634))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111011" => if(ecg(636) > ecg(635))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(636))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(635)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(636) < ecg(635))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(635))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(636)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(635))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111100" => if(ecg(637) > ecg(636))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(637))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(636)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(637) < ecg(636))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(636))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(637)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(636))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111101" => if(ecg(638) > ecg(637))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(638))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(637)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(638) < ecg(637))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(637))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(638)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(637))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111110" => if(ecg(639) > ecg(638))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(639))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(638)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        elsif(ecg(639) < ecg(638))then
                          if((conv_integer(v_counter) >= (conv_integer(v_distance_c) - conv_integer(ecg(638))))
                             and (conv_integer(v_counter) <= (conv_integer(v_distance_c) - conv_integer(ecg(639)))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        else
                          if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(638))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                          else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                          end if;
                        end if;

 when "1001111111" => if(conv_integer(v_counter) = (conv_integer(v_distance_c) - conv_integer(ecg(639))))then
                                                   red   <= "111";
                                                   green <= "100";
                                                   blue  <=  "00";
                        else
                                                   red   <= "000";
                                                   green <= "000";
                                                   blue  <=  "00";
                        end if;
                                           
 when others =>         red   <= "000";
                        green <= "000";
                        blue  <=  "00";
 end case;

 end if;

 end process image_p;

end Behavioral;