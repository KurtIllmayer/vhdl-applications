----------------------------------------------------------------------------------
--
-- Company:         Bulme Graz Goesting
-- Engineer:        Kurt Illmayer
-- 
-- Creation Date:   18:25:33 02/15/2019
-- Design Name:     test10
-- Module Name:     test10 - Behavioral
-- File Name:       C:/Digital_Designs/SCHILF_VHDL/VHDL_Applications/count_ones/test10.vhd
-- Project Name:    VHDL Applications
-- Target Devices:  XC3S100E
-- Tool versions:   ISE Webpack 14.7
-- Description:     VHDL Basic Designs
--
-- Revision 0.1 -   File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity test10 is
    Port ( a_i : in  STD_ULOGIC;
           b_i : in  STD_ULOGIC;
           c_o : out  STD_ULOGIC);
end test10;

architecture Behavioral of test10 is

begin


end Behavioral;
